module VNLP_TB;
	
	wire [26:0] Result;
	wire [7:0] Len;
	wire Done;
	wire [8:0] A1;
	wire [8:0] A2;
	wire [9:0] D1;
	wire [9:0] D2;
	reg Start;
	reg Reset;
	reg Clk;
	

	VNLP underTest(
		.Result(Result),
		.Len(Len),
		.Done(Done),
		.Start(Start),
		.Reset(Reset),
		.Clk(Clk));

	assign A1= underTest.MemAdd1;
	assign A2= underTest.MemAdd2;
	assign D1= underTest.MemData1;
	assign D2= underTest.MemData2;

	reg [9:0] k;
	initial begin: Flush_Memory
		#2 for (k= 0; k < 512; k=k+1) underTest.M.Data[k]= 0;
	end
 
	initial begin: Initialize_Values
		Clk= 0;
		#7
		Start= 0;
		Reset= 1;
		#1
		Reset= 0;
		Start= 1;
		#7
		Start= 0;
	end

	initial begin: Load_List
		#5
		underTest.M.Data[0]= 10'b0000110001;
		underTest.M.Data[1]= 10'b0000100010;
		underTest.M.Data[2]= 10'b1111011111;
		underTest.M.Data[3]= 10'b0000010111;
		underTest.M.Data[5]= 10'b0000010001;
		underTest.M.Data[6]= 10'b0000101000;
		underTest.M.Data[7]= 10'b0000010011;
		underTest.M.Data[8]= 10'b0001100110;
		underTest.M.Data[11]= 10'b0000010110;
		underTest.M.Data[12]= 10'b0000010010;
		underTest.M.Data[13]= 10'b0000011001;
		underTest.M.Data[14]= 10'b1110100011;
		underTest.M.Data[17]= 10'b0000001011;
		underTest.M.Data[18]= 10'b0000000110;
		underTest.M.Data[19]= 10'b0000001000;
		underTest.M.Data[20]= 10'b0001011010;
		underTest.M.Data[22]= 10'b0000100001;
		underTest.M.Data[23]= 10'b0000001100;
		underTest.M.Data[24]= 10'b0000011111;
		underTest.M.Data[25]= 10'b0000100000;
		underTest.M.Data[28]= 10'b0001100110;
		underTest.M.Data[29]= 10'b0011110000;
		underTest.M.Data[30]= 10'b0000101111;
		underTest.M.Data[31]= 10'b1111110101;
		underTest.M.Data[33]= 10'b0000000000;
		underTest.M.Data[34]= 10'b0000010111;
		underTest.M.Data[35]= 10'b0000011001;
		underTest.M.Data[36]= 10'b0001011000;
		underTest.M.Data[39]= 10'b0000000101;
		underTest.M.Data[40]= 10'b0000110010;
		underTest.M.Data[41]= 10'b0000111000;
		underTest.M.Data[42]= 10'b0000110000;
		underTest.M.Data[44]= 10'b0000111000;
		underTest.M.Data[45]= 10'b0001011000;
		underTest.M.Data[46]= 10'b0001110000;
		underTest.M.Data[47]= 10'b0001000101;
		underTest.M.Data[49]= 10'b0000100111;
		underTest.M.Data[50]= 10'b0000000001;
		underTest.M.Data[51]= 10'b0001100101;
		underTest.M.Data[52]= 10'b0000111111;
	end

	always begin
		#10 Clk= ~Clk;
	end

endmodule

module VNLP_TB2;
	
	wire [26:0] Result;
	wire [7:0] Len;
	wire Done;
	wire [8:0] A1;
	wire [8:0] A2;
	wire [9:0] D1;
	wire [9:0] D2;
	reg Start;
	reg Reset;
	reg Clk;
	
	VNLP underTest(
		.Result(Result),
		.Len(Len),
		.Done(Done),
		.Start(Start),
		.Reset(Reset),
		.Clk(Clk));

	assign A1= underTest.MemAdd1;
	assign A2= underTest.MemAdd2;
	assign D1= underTest.MemData1;
	assign D2= underTest.MemData2;


	reg [9:0] k;
	initial begin: Flush_Memory
		#2 for (k= 0; k < 512; k=k+1) underTest.M.Data[k]= 0;
	end
 
	initial begin: Initialize_Values
		Clk= 0;
		#7
		Start= 0;
		Reset= 1;
		#1
		Reset= 0;
		Start= 1;
		#7
		Start= 0;
	end

	initial begin: Load_List
		#5
		underTest.M.Data[0]= 10'd4;
		underTest.M.Data[1]= 10'd509;
		underTest.M.Data[2]= -10'sd512;
		underTest.M.Data[3]= -10'sd512;
		underTest.M.Data[4]= 10'd8;
		underTest.M.Data[5]= 10'd1;
		underTest.M.Data[6]= -10'sd512;
		underTest.M.Data[7]= -10'sd512;
		underTest.M.Data[8]= 10'd12;
		underTest.M.Data[9]= 10'd5;
		underTest.M.Data[10]= -10'sd512;
		underTest.M.Data[11]= -10'sd512;
		underTest.M.Data[12]= 10'd16;
		underTest.M.Data[13]= 10'd9;
		underTest.M.Data[14]= -10'sd512;
		underTest.M.Data[15]= -10'sd512;
		underTest.M.Data[16]= 10'd20;
		underTest.M.Data[17]= 10'd13;
		underTest.M.Data[18]= -10'sd512;
		underTest.M.Data[19]= -10'sd512;
		underTest.M.Data[20]= 10'd24;
		underTest.M.Data[21]= 10'd17;
		underTest.M.Data[22]= -10'sd512;
		underTest.M.Data[23]= -10'sd512;
		underTest.M.Data[24]= 10'd28;
		underTest.M.Data[25]= 10'd21;
		underTest.M.Data[26]= -10'sd512;
		underTest.M.Data[27]= -10'sd512;
		underTest.M.Data[28]= 10'd32;
		underTest.M.Data[29]= 10'd25;
		underTest.M.Data[30]= -10'sd512;
		underTest.M.Data[31]= -10'sd512;
		underTest.M.Data[32]= 10'd36;
		underTest.M.Data[33]= 10'd29;
		underTest.M.Data[34]= -10'sd512;
		underTest.M.Data[35]= -10'sd512;
		underTest.M.Data[36]= 10'd40;
		underTest.M.Data[37]= 10'd33;
		underTest.M.Data[38]= -10'sd512;
		underTest.M.Data[39]= -10'sd512;
		underTest.M.Data[40]= 10'd44;
		underTest.M.Data[41]= 10'd37;
		underTest.M.Data[42]= -10'sd512;
		underTest.M.Data[43]= -10'sd512;
		underTest.M.Data[44]= 10'd48;
		underTest.M.Data[45]= 10'd41;
		underTest.M.Data[46]= -10'sd512;
		underTest.M.Data[47]= -10'sd512;
		underTest.M.Data[48]= 10'd52;
		underTest.M.Data[49]= 10'd45;
		underTest.M.Data[50]= -10'sd512;
		underTest.M.Data[51]= -10'sd512;
		underTest.M.Data[52]= 10'd56;
		underTest.M.Data[53]= 10'd49;
		underTest.M.Data[54]= -10'sd512;
		underTest.M.Data[55]= -10'sd512;
		underTest.M.Data[56]= 10'd60;
		underTest.M.Data[57]= 10'd53;
		underTest.M.Data[58]= -10'sd512;
		underTest.M.Data[59]= -10'sd512;
		underTest.M.Data[60]= 10'd64;
		underTest.M.Data[61]= 10'd57;
		underTest.M.Data[62]= -10'sd512;
		underTest.M.Data[63]= -10'sd512;
		underTest.M.Data[64]= 10'd68;
		underTest.M.Data[65]= 10'd61;
		underTest.M.Data[66]= -10'sd512;
		underTest.M.Data[67]= -10'sd512;
		underTest.M.Data[68]= 10'd72;
		underTest.M.Data[69]= 10'd65;
		underTest.M.Data[70]= -10'sd512;
		underTest.M.Data[71]= -10'sd512;
		underTest.M.Data[72]= 10'd76;
		underTest.M.Data[73]= 10'd69;
		underTest.M.Data[74]= -10'sd512;
		underTest.M.Data[75]= -10'sd512;
		underTest.M.Data[76]= 10'd80;
		underTest.M.Data[77]= 10'd73;
		underTest.M.Data[78]= -10'sd512;
		underTest.M.Data[79]= -10'sd512;
		underTest.M.Data[80]= 10'd84;
		underTest.M.Data[81]= 10'd77;
		underTest.M.Data[82]= -10'sd512;
		underTest.M.Data[83]= -10'sd512;
		underTest.M.Data[84]= 10'd88;
		underTest.M.Data[85]= 10'd81;
		underTest.M.Data[86]= -10'sd512;
		underTest.M.Data[87]= -10'sd512;
		underTest.M.Data[88]= 10'd92;
		underTest.M.Data[89]= 10'd85;
		underTest.M.Data[90]= -10'sd512;
		underTest.M.Data[91]= -10'sd512;
		underTest.M.Data[92]= 10'd96;
		underTest.M.Data[93]= 10'd89;
		underTest.M.Data[94]= -10'sd512;
		underTest.M.Data[95]= -10'sd512;
		underTest.M.Data[96]= 10'd100;
		underTest.M.Data[97]= 10'd93;
		underTest.M.Data[98]= -10'sd512;
		underTest.M.Data[99]= -10'sd512;
		underTest.M.Data[100]= 10'd104;
		underTest.M.Data[101]= 10'd97;
		underTest.M.Data[102]= -10'sd512;
		underTest.M.Data[103]= -10'sd512;
		underTest.M.Data[104]= 10'd108;
		underTest.M.Data[105]= 10'd101;
		underTest.M.Data[106]= -10'sd512;
		underTest.M.Data[107]= -10'sd512;
		underTest.M.Data[108]= 10'd112;
		underTest.M.Data[109]= 10'd105;
		underTest.M.Data[110]= -10'sd512;
		underTest.M.Data[111]= -10'sd512;
		underTest.M.Data[112]= 10'd116;
		underTest.M.Data[113]= 10'd109;
		underTest.M.Data[114]= -10'sd512;
		underTest.M.Data[115]= -10'sd512;
		underTest.M.Data[116]= 10'd120;
		underTest.M.Data[117]= 10'd113;
		underTest.M.Data[118]= -10'sd512;
		underTest.M.Data[119]= -10'sd512;
		underTest.M.Data[120]= 10'd124;
		underTest.M.Data[121]= 10'd117;
		underTest.M.Data[122]= -10'sd512;
		underTest.M.Data[123]= -10'sd512;
		underTest.M.Data[124]= 10'd128;
		underTest.M.Data[125]= 10'd121;
		underTest.M.Data[126]= -10'sd512;
		underTest.M.Data[127]= -10'sd512;
		underTest.M.Data[128]= 10'd132;
		underTest.M.Data[129]= 10'd125;
		underTest.M.Data[130]= -10'sd512;
		underTest.M.Data[131]= -10'sd512;
		underTest.M.Data[132]= 10'd136;
		underTest.M.Data[133]= 10'd129;
		underTest.M.Data[134]= -10'sd512;
		underTest.M.Data[135]= -10'sd512;
		underTest.M.Data[136]= 10'd140;
		underTest.M.Data[137]= 10'd133;
		underTest.M.Data[138]= -10'sd512;
		underTest.M.Data[139]= -10'sd512;
		underTest.M.Data[140]= 10'd144;
		underTest.M.Data[141]= 10'd137;
		underTest.M.Data[142]= -10'sd512;
		underTest.M.Data[143]= -10'sd512;
		underTest.M.Data[144]= 10'd148;
		underTest.M.Data[145]= 10'd141;
		underTest.M.Data[146]= -10'sd512;
		underTest.M.Data[147]= -10'sd512;
		underTest.M.Data[148]= 10'd152;
		underTest.M.Data[149]= 10'd145;
		underTest.M.Data[150]= -10'sd512;
		underTest.M.Data[151]= -10'sd512;
		underTest.M.Data[152]= 10'd156;
		underTest.M.Data[153]= 10'd149;
		underTest.M.Data[154]= -10'sd512;
		underTest.M.Data[155]= -10'sd512;
		underTest.M.Data[156]= 10'd160;
		underTest.M.Data[157]= 10'd153;
		underTest.M.Data[158]= -10'sd512;
		underTest.M.Data[159]= -10'sd512;
		underTest.M.Data[160]= 10'd164;
		underTest.M.Data[161]= 10'd157;
		underTest.M.Data[162]= -10'sd512;
		underTest.M.Data[163]= -10'sd512;
		underTest.M.Data[164]= 10'd168;
		underTest.M.Data[165]= 10'd161;
		underTest.M.Data[166]= -10'sd512;
		underTest.M.Data[167]= -10'sd512;
		underTest.M.Data[168]= 10'd172;
		underTest.M.Data[169]= 10'd165;
		underTest.M.Data[170]= -10'sd512;
		underTest.M.Data[171]= -10'sd512;
		underTest.M.Data[172]= 10'd176;
		underTest.M.Data[173]= 10'd169;
		underTest.M.Data[174]= -10'sd512;
		underTest.M.Data[175]= -10'sd512;
		underTest.M.Data[176]= 10'd180;
		underTest.M.Data[177]= 10'd173;
		underTest.M.Data[178]= -10'sd512;
		underTest.M.Data[179]= -10'sd512;
		underTest.M.Data[180]= 10'd184;
		underTest.M.Data[181]= 10'd177;
		underTest.M.Data[182]= -10'sd512;
		underTest.M.Data[183]= -10'sd512;
		underTest.M.Data[184]= 10'd188;
		underTest.M.Data[185]= 10'd181;
		underTest.M.Data[186]= -10'sd512;
		underTest.M.Data[187]= -10'sd512;
		underTest.M.Data[188]= 10'd192;
		underTest.M.Data[189]= 10'd185;
		underTest.M.Data[190]= -10'sd512;
		underTest.M.Data[191]= -10'sd512;
		underTest.M.Data[192]= 10'd196;
		underTest.M.Data[193]= 10'd189;
		underTest.M.Data[194]= -10'sd512;
		underTest.M.Data[195]= -10'sd512;
		underTest.M.Data[196]= 10'd200;
		underTest.M.Data[197]= 10'd193;
		underTest.M.Data[198]= -10'sd512;
		underTest.M.Data[199]= -10'sd512;
		underTest.M.Data[200]= 10'd204;
		underTest.M.Data[201]= 10'd197;
		underTest.M.Data[202]= -10'sd512;
		underTest.M.Data[203]= -10'sd512;
		underTest.M.Data[204]= 10'd208;
		underTest.M.Data[205]= 10'd201;
		underTest.M.Data[206]= -10'sd512;
		underTest.M.Data[207]= -10'sd512;
		underTest.M.Data[208]= 10'd212;
		underTest.M.Data[209]= 10'd205;
		underTest.M.Data[210]= -10'sd512;
		underTest.M.Data[211]= -10'sd512;
		underTest.M.Data[212]= 10'd216;
		underTest.M.Data[213]= 10'd209;
		underTest.M.Data[214]= -10'sd512;
		underTest.M.Data[215]= -10'sd512;
		underTest.M.Data[216]= 10'd220;
		underTest.M.Data[217]= 10'd213;
		underTest.M.Data[218]= -10'sd512;
		underTest.M.Data[219]= -10'sd512;
		underTest.M.Data[220]= 10'd224;
		underTest.M.Data[221]= 10'd217;
		underTest.M.Data[222]= -10'sd512;
		underTest.M.Data[223]= -10'sd512;
		underTest.M.Data[224]= 10'd228;
		underTest.M.Data[225]= 10'd221;
		underTest.M.Data[226]= -10'sd512;
		underTest.M.Data[227]= -10'sd512;
		underTest.M.Data[228]= 10'd232;
		underTest.M.Data[229]= 10'd225;
		underTest.M.Data[230]= -10'sd512;
		underTest.M.Data[231]= -10'sd512;
		underTest.M.Data[232]= 10'd236;
		underTest.M.Data[233]= 10'd229;
		underTest.M.Data[234]= -10'sd512;
		underTest.M.Data[235]= -10'sd512;
		underTest.M.Data[236]= 10'd240;
		underTest.M.Data[237]= 10'd233;
		underTest.M.Data[238]= -10'sd512;
		underTest.M.Data[239]= -10'sd512;
		underTest.M.Data[240]= 10'd244;
		underTest.M.Data[241]= 10'd237;
		underTest.M.Data[242]= -10'sd512;
		underTest.M.Data[243]= -10'sd512;
		underTest.M.Data[244]= 10'd248;
		underTest.M.Data[245]= 10'd241;
		underTest.M.Data[246]= -10'sd512;
		underTest.M.Data[247]= -10'sd512;
		underTest.M.Data[248]= 10'd252;
		underTest.M.Data[249]= 10'd245;
		underTest.M.Data[250]= -10'sd512;
		underTest.M.Data[251]= -10'sd512;
		underTest.M.Data[252]= 10'd256;
		underTest.M.Data[253]= 10'd249;
		underTest.M.Data[254]= -10'sd512;
		underTest.M.Data[255]= -10'sd512;
		underTest.M.Data[256]= 10'd260;
		underTest.M.Data[257]= 10'd253;
		underTest.M.Data[258]= -10'sd512;
		underTest.M.Data[259]= -10'sd512;
		underTest.M.Data[260]= 10'd264;
		underTest.M.Data[261]= 10'd257;
		underTest.M.Data[262]= -10'sd512;
		underTest.M.Data[263]= -10'sd512;
		underTest.M.Data[264]= 10'd268;
		underTest.M.Data[265]= 10'd261;
		underTest.M.Data[266]= -10'sd512;
		underTest.M.Data[267]= -10'sd512;
		underTest.M.Data[268]= 10'd272;
		underTest.M.Data[269]= 10'd265;
		underTest.M.Data[270]= -10'sd512;
		underTest.M.Data[271]= -10'sd512;
		underTest.M.Data[272]= 10'd276;
		underTest.M.Data[273]= 10'd269;
		underTest.M.Data[274]= -10'sd512;
		underTest.M.Data[275]= -10'sd512;
		underTest.M.Data[276]= 10'd280;
		underTest.M.Data[277]= 10'd273;
		underTest.M.Data[278]= -10'sd512;
		underTest.M.Data[279]= -10'sd512;
		underTest.M.Data[280]= 10'd284;
		underTest.M.Data[281]= 10'd277;
		underTest.M.Data[282]= -10'sd512;
		underTest.M.Data[283]= -10'sd512;
		underTest.M.Data[284]= 10'd288;
		underTest.M.Data[285]= 10'd281;
		underTest.M.Data[286]= -10'sd512;
		underTest.M.Data[287]= -10'sd512;
		underTest.M.Data[288]= 10'd292;
		underTest.M.Data[289]= 10'd285;
		underTest.M.Data[290]= -10'sd512;
		underTest.M.Data[291]= -10'sd512;
		underTest.M.Data[292]= 10'd296;
		underTest.M.Data[293]= 10'd289;
		underTest.M.Data[294]= -10'sd512;
		underTest.M.Data[295]= -10'sd512;
		underTest.M.Data[296]= 10'd300;
		underTest.M.Data[297]= 10'd293;
		underTest.M.Data[298]= -10'sd512;
		underTest.M.Data[299]= -10'sd512;
		underTest.M.Data[300]= 10'd304;
		underTest.M.Data[301]= 10'd297;
		underTest.M.Data[302]= -10'sd512;
		underTest.M.Data[303]= -10'sd512;
		underTest.M.Data[304]= 10'd308;
		underTest.M.Data[305]= 10'd301;
		underTest.M.Data[306]= -10'sd512;
		underTest.M.Data[307]= -10'sd512;
		underTest.M.Data[308]= 10'd312;
		underTest.M.Data[309]= 10'd305;
		underTest.M.Data[310]= -10'sd512;
		underTest.M.Data[311]= -10'sd512;
		underTest.M.Data[312]= 10'd316;
		underTest.M.Data[313]= 10'd309;
		underTest.M.Data[314]= -10'sd512;
		underTest.M.Data[315]= -10'sd512;
		underTest.M.Data[316]= 10'd320;
		underTest.M.Data[317]= 10'd313;
		underTest.M.Data[318]= -10'sd512;
		underTest.M.Data[319]= -10'sd512;
		underTest.M.Data[320]= 10'd324;
		underTest.M.Data[321]= 10'd317;
		underTest.M.Data[322]= -10'sd512;
		underTest.M.Data[323]= -10'sd512;
		underTest.M.Data[324]= 10'd328;
		underTest.M.Data[325]= 10'd321;
		underTest.M.Data[326]= -10'sd512;
		underTest.M.Data[327]= -10'sd512;
		underTest.M.Data[328]= 10'd332;
		underTest.M.Data[329]= 10'd325;
		underTest.M.Data[330]= -10'sd512;
		underTest.M.Data[331]= -10'sd512;
		underTest.M.Data[332]= 10'd336;
		underTest.M.Data[333]= 10'd329;
		underTest.M.Data[334]= -10'sd512;
		underTest.M.Data[335]= -10'sd512;
		underTest.M.Data[336]= 10'd340;
		underTest.M.Data[337]= 10'd333;
		underTest.M.Data[338]= -10'sd512;
		underTest.M.Data[339]= -10'sd512;
		underTest.M.Data[340]= 10'd344;
		underTest.M.Data[341]= 10'd337;
		underTest.M.Data[342]= -10'sd512;
		underTest.M.Data[343]= -10'sd512;
		underTest.M.Data[344]= 10'd348;
		underTest.M.Data[345]= 10'd341;
		underTest.M.Data[346]= -10'sd512;
		underTest.M.Data[347]= -10'sd512;
		underTest.M.Data[348]= 10'd352;
		underTest.M.Data[349]= 10'd345;
		underTest.M.Data[350]= -10'sd512;
		underTest.M.Data[351]= -10'sd512;
		underTest.M.Data[352]= 10'd356;
		underTest.M.Data[353]= 10'd349;
		underTest.M.Data[354]= -10'sd512;
		underTest.M.Data[355]= -10'sd512;
		underTest.M.Data[356]= 10'd360;
		underTest.M.Data[357]= 10'd353;
		underTest.M.Data[358]= -10'sd512;
		underTest.M.Data[359]= -10'sd512;
		underTest.M.Data[360]= 10'd364;
		underTest.M.Data[361]= 10'd357;
		underTest.M.Data[362]= -10'sd512;
		underTest.M.Data[363]= -10'sd512;
		underTest.M.Data[364]= 10'd368;
		underTest.M.Data[365]= 10'd361;
		underTest.M.Data[366]= -10'sd512;
		underTest.M.Data[367]= -10'sd512;
		underTest.M.Data[368]= 10'd372;
		underTest.M.Data[369]= 10'd365;
		underTest.M.Data[370]= -10'sd512;
		underTest.M.Data[371]= -10'sd512;
		underTest.M.Data[372]= 10'd376;
		underTest.M.Data[373]= 10'd369;
		underTest.M.Data[374]= -10'sd512;
		underTest.M.Data[375]= -10'sd512;
		underTest.M.Data[376]= 10'd380;
		underTest.M.Data[377]= 10'd373;
		underTest.M.Data[378]= -10'sd512;
		underTest.M.Data[379]= -10'sd512;
		underTest.M.Data[380]= 10'd384;
		underTest.M.Data[381]= 10'd377;
		underTest.M.Data[382]= -10'sd512;
		underTest.M.Data[383]= -10'sd512;
		underTest.M.Data[384]= 10'd388;
		underTest.M.Data[385]= 10'd381;
		underTest.M.Data[386]= -10'sd512;
		underTest.M.Data[387]= -10'sd512;
		underTest.M.Data[388]= 10'd392;
		underTest.M.Data[389]= 10'd385;
		underTest.M.Data[390]= -10'sd512;
		underTest.M.Data[391]= -10'sd512;
		underTest.M.Data[392]= 10'd396;
		underTest.M.Data[393]= 10'd389;
		underTest.M.Data[394]= -10'sd512;
		underTest.M.Data[395]= -10'sd512;
		underTest.M.Data[396]= 10'd400;
		underTest.M.Data[397]= 10'd393;
		underTest.M.Data[398]= -10'sd512;
		underTest.M.Data[399]= -10'sd512;
		underTest.M.Data[400]= 10'd404;
		underTest.M.Data[401]= 10'd397;
		underTest.M.Data[402]= -10'sd512;
		underTest.M.Data[403]= -10'sd512;
		underTest.M.Data[404]= 10'd408;
		underTest.M.Data[405]= 10'd401;
		underTest.M.Data[406]= -10'sd512;
		underTest.M.Data[407]= -10'sd512;
		underTest.M.Data[408]= 10'd412;
		underTest.M.Data[409]= 10'd405;
		underTest.M.Data[410]= -10'sd512;
		underTest.M.Data[411]= -10'sd512;
		underTest.M.Data[412]= 10'd416;
		underTest.M.Data[413]= 10'd409;
		underTest.M.Data[414]= -10'sd512;
		underTest.M.Data[415]= -10'sd512;
		underTest.M.Data[416]= 10'd420;
		underTest.M.Data[417]= 10'd413;
		underTest.M.Data[418]= -10'sd512;
		underTest.M.Data[419]= -10'sd512;
		underTest.M.Data[420]= 10'd424;
		underTest.M.Data[421]= 10'd417;
		underTest.M.Data[422]= -10'sd512;
		underTest.M.Data[423]= -10'sd512;
		underTest.M.Data[424]= 10'd428;
		underTest.M.Data[425]= 10'd421;
		underTest.M.Data[426]= -10'sd512;
		underTest.M.Data[427]= -10'sd512;
		underTest.M.Data[428]= 10'd432;
		underTest.M.Data[429]= 10'd425;
		underTest.M.Data[430]= -10'sd512;
		underTest.M.Data[431]= -10'sd512;
		underTest.M.Data[432]= 10'd436;
		underTest.M.Data[433]= 10'd429;
		underTest.M.Data[434]= -10'sd512;
		underTest.M.Data[435]= -10'sd512;
		underTest.M.Data[436]= 10'd440;
		underTest.M.Data[437]= 10'd433;
		underTest.M.Data[438]= -10'sd512;
		underTest.M.Data[439]= -10'sd512;
		underTest.M.Data[440]= 10'd444;
		underTest.M.Data[441]= 10'd437;
		underTest.M.Data[442]= -10'sd512;
		underTest.M.Data[443]= -10'sd512;
		underTest.M.Data[444]= 10'd448;
		underTest.M.Data[445]= 10'd441;
		underTest.M.Data[446]= -10'sd512;
		underTest.M.Data[447]= -10'sd512;
		underTest.M.Data[448]= 10'd452;
		underTest.M.Data[449]= 10'd445;
		underTest.M.Data[450]= -10'sd512;
		underTest.M.Data[451]= -10'sd512;
		underTest.M.Data[452]= 10'd456;
		underTest.M.Data[453]= 10'd449;
		underTest.M.Data[454]= -10'sd512;
		underTest.M.Data[455]= -10'sd512;
		underTest.M.Data[456]= 10'd460;
		underTest.M.Data[457]= 10'd453;
		underTest.M.Data[458]= -10'sd512;
		underTest.M.Data[459]= -10'sd512;
		underTest.M.Data[460]= 10'd464;
		underTest.M.Data[461]= 10'd457;
		underTest.M.Data[462]= -10'sd512;
		underTest.M.Data[463]= -10'sd512;
		underTest.M.Data[464]= 10'd468;
		underTest.M.Data[465]= 10'd461;
		underTest.M.Data[466]= -10'sd512;
		underTest.M.Data[467]= -10'sd512;
		underTest.M.Data[468]= 10'd472;
		underTest.M.Data[469]= 10'd465;
		underTest.M.Data[470]= -10'sd512;
		underTest.M.Data[471]= -10'sd512;
		underTest.M.Data[472]= 10'd476;
		underTest.M.Data[473]= 10'd469;
		underTest.M.Data[474]= -10'sd512;
		underTest.M.Data[475]= -10'sd512;
		underTest.M.Data[476]= 10'd480;
		underTest.M.Data[477]= 10'd473;
		underTest.M.Data[478]= -10'sd512;
		underTest.M.Data[479]= -10'sd512;
		underTest.M.Data[480]= 10'd484;
		underTest.M.Data[481]= 10'd477;
		underTest.M.Data[482]= -10'sd512;
		underTest.M.Data[483]= -10'sd512;
		underTest.M.Data[484]= 10'd488;
		underTest.M.Data[485]= 10'd481;
		underTest.M.Data[486]= -10'sd512;
		underTest.M.Data[487]= -10'sd512;
		underTest.M.Data[488]= 10'd492;
		underTest.M.Data[489]= 10'd485;
		underTest.M.Data[490]= -10'sd512;
		underTest.M.Data[491]= -10'sd512;
		underTest.M.Data[492]= 10'd496;
		underTest.M.Data[493]= 10'd489;
		underTest.M.Data[494]= -10'sd512;
		underTest.M.Data[495]= -10'sd512;
		underTest.M.Data[496]= 10'd500;
		underTest.M.Data[497]= 10'd493;
		underTest.M.Data[498]= -10'sd512;
		underTest.M.Data[499]= -10'sd512;
		underTest.M.Data[500]= 10'd504;
		underTest.M.Data[501]= 10'd497;
		underTest.M.Data[502]= -10'sd512;
		underTest.M.Data[503]= -10'sd512;
		underTest.M.Data[504]= 10'd508;
		underTest.M.Data[505]= 10'd501;
		underTest.M.Data[506]= -10'sd512;
		underTest.M.Data[507]= -10'sd512;
		underTest.M.Data[508]= 10'd0;
		underTest.M.Data[509]= 10'd505;
		underTest.M.Data[510]= -10'sd512;
		underTest.M.Data[511]= -10'sd512;
	end

	always begin
		#10 Clk= ~Clk;
	end

endmodule